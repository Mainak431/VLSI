*** SPICE deck for cell inverter{ic} from library INV
*** Created on Thu Jul 21, 2016 21:55:51
*** Last revised on Fri Jul 22, 2016 00:30:07
*** Written on Fri Jul 22, 2016 00:32:01 by Electric VLSI Design System, 
*version 9.04
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.OPTIONS NOMOD DEFL=3UM DEFW=3UM DEFAD=70P DEFAS=70P LIMPTS=1000
+ITL5=0 RELTOL=0.01 ABSTOL=500PA VNTOL=500UV LVLTIM=2
+LVLCOD=1
.MODEL N NMOS LEVEL=1
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL P PMOS LEVEL=1
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2

*** TOP LEVEL CELL: INV:inverter{ic}

* Spice Code nodes in cell cell 'INV:inverter{ic}'
vdd vdd 0 DC 5
vin in 0 DC 0
.dc vin 0 5 1m
.include C:\Users\Mainak\Desktop\vlsi\32nm_hp.txt
.END
